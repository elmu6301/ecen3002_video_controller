/*
    ECEN 3002
    Video Project: Reset Module
    Elena Murray

*/

// module reset(
    
// ); 

// endmodule